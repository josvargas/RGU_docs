/**********************************************************************************
Theia, Ray Cast Programable graphic Processing Unit.
Copyright (C) 2014  Diego Valverde (diego.valverde.g@gmail.com)

This program is free software; you can redistribute it and/or
modify it under the terms of the GNU General Public License
as published by the Free Software Foundation; either version 2
of the License, or (at your option) any later version.

This program is distributed in the hope that it will be useful,
but WITHOUT ANY WARRANTY; without even the implied warranty of
MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
GNU General Public License for more details.

You should have received a copy of the GNU General Public License
along with this program; if not, write to the Free Software
Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.

***********************************************************************************/
`timescale 1ns / 1ps

`include "Definitions.v"

module SimpleOperationTestBench;

	// Inputs
	reg iClock;
	reg iReset;
	reg iEnable;
	reg iUartSelected;
	reg iUartWrite;
	reg [7:0] iUartAddr;
	reg [`GPU_WORD-1:0] iUartData;

	// Outputs
	wire oFifoPush;
	wire [`GPU_WORD-1:0] oFifoData;
	wire [`GPU_WORD-1:0] oUartData;	

	always
	begin
		repeat(3000) begin
			#`GLOBAL_CLOCK_CYCLE iClock = ~iClock;
		end
		$finish;
	end

	// Instantiate the Unit Under Test (UUT)
	RayGenerationUnit RGU (
		.iClock(iClock),
		.iReset(iReset),
	 	.iEnable(iEnable),
		.oFifoPush(oFifoPush),
		.oFifoData(oFifoData),
		.iUartSelected(iUartSelected),
		.iUartWrite(iUartWrite),
		.iUartAddr(iUartAddr),
		.iUartData(iUartData),
		.oUartData(oUartData)
	);

	reg [`RGU_RANDOM_SIZE-1:0] random;

	`include "driver.v"
	`include "checker_3.v"

	parameter ITERATIONS = 3000;
	integer log;

	initial begin

		$dumpfile("rgu.vcd");
		$dumpvars;

		log = $fopen("tb_3.log");

		// Initialize Inputs
		iClock = 0;
		iReset = 0;
		iEnable = 1;
		// Wait 100 ns for global reset to finish
		#100;
		iReset = 1;
		RGU.INSTRUCTION_RAM.Ram[0] = {`CONTINUE, `NOBREAK, 1'b0,`RGU_SQRT ,5'd7,5'd1,5'd1};
		#(50*`GLOBAL_CLOCK_PERIOD)
		iReset = 0;
		
		//random = $random;
		RGU.DATA_RAM.Ram[0] = 32'h0;		
		//RGU.DATA_RAM.Ram[1] = 32'h40000;
		RGU.DATA_RAM.Ram[1] = {11'b0,4'b0010,17'b0};			
		RGU.DATA_RAM.Ram[2] = 32'h60000;
		RGU.DATA_RAM.Ram[3] = 32'h40000;
		RGU.DATA_RAM.Ram[4] = 32'h20000;

		RGU.INSTRUCTION_RAM.Ram[0] = {`CONTINUE, `NOBREAK, 1'b0,`RGU_SQRT ,5'd7,5'd1,5'd1};
		RGU.INSTRUCTION_RAM.Ram[1] = {`CONTINUE, `NOBREAK, 1'b0,`RGU_MUL  ,5'd8,5'd7,5'd7};
		RGU.INSTRUCTION_RAM.Ram[2] = {`CONTINUE, `NOBREAK, 1'b0,`RGU_MUL  ,5'd9,5'd1,5'd8};
		RGU.INSTRUCTION_RAM.Ram[3] = {`CONTINUE, `NOBREAK, 1'b0,`RGU_SUB  ,5'd10,5'd2,5'd9};
		RGU.INSTRUCTION_RAM.Ram[4] = {`CONTINUE, `NOBREAK, 1'b0,`RGU_MUL  ,5'd11,5'd10,5'd7};
		RGU.INSTRUCTION_RAM.Ram[5] = {`CONTINUE, `NOBREAK, 1'b0,`RGU_DIV  ,5'd12,5'd11,5'd3};
		RGU.INSTRUCTION_RAM.Ram[6] = {`CONTINUE, `NOBREAK, 1'b0,`RGU_MUL  ,5'd8,5'd12,5'd12};
		RGU.INSTRUCTION_RAM.Ram[7] = {`CONTINUE, `NOBREAK, 1'b0,`RGU_MUL  ,5'd9,5'd1,5'd8};
		RGU.INSTRUCTION_RAM.Ram[8] = {`CONTINUE, `NOBREAK, 1'b0,`RGU_SUB  ,5'd10,5'd2,5'd9};
		RGU.INSTRUCTION_RAM.Ram[9] = {`CONTINUE, `NOBREAK, 1'b0,`RGU_MUL  ,5'd11,5'd10,5'd12};
		RGU.INSTRUCTION_RAM.Ram[10] = {`CONTINUE, `NOBREAK, 1'b0,`RGU_DIV  ,5'd13,5'd11,5'd3};
		RGU.INSTRUCTION_RAM.Ram[11] = {`CONTINUE, `NOBREAK, 1'b0,`RGU_MUL  ,5'd8,5'd13,5'd13};
		RGU.INSTRUCTION_RAM.Ram[12] = {`CONTINUE, `NOBREAK, 1'b0,`RGU_MUL  ,5'd9,5'd1,5'd8};
		RGU.INSTRUCTION_RAM.Ram[13] = {`CONTINUE, `NOBREAK, 1'b0,`RGU_SUB  ,5'd10,5'd2,5'd9};
		RGU.INSTRUCTION_RAM.Ram[14] = {`CONTINUE, `NOBREAK, 1'b0,`RGU_MUL  ,5'd11,5'd10,5'd13};
		RGU.INSTRUCTION_RAM.Ram[15] = {`CONTINUE, `NOBREAK, 1'b0,`RGU_DIV  ,5'd12,5'd11,5'd3};				
		RGU.INSTRUCTION_RAM.Ram[16] = {`CONTINUE, `NOBREAK, 1'b0,`RGU_PUSH  ,5'd0,5'd12,5'd0};

		fork
			drv_random(ITERATIONS);
			drv_ram(ITERATIONS);
			checker(ITERATIONS);
		join

		$fclose(log);
		//#200 $finish;

		//$display("%x",RGU.DATA_RAM.Ram[1]);

	end
      
endmodule 
